package Stage1;

	(*synthesize*)
	module mkStage1(Empty);	
		Mem instMem <- mkMem(INST_CACHE_SIZE);
	
		
	
	endmodule: mkStage1


endpackage
