package Stage5;

	`include "Constants.defines"
	import Utils::*;
	import PipeRegs::*;
	
	module mkStage5 #(MemWb memWb) (Empty);
	
	endmodule: mkStage5
endpackage
