package DataTypes;

	typedef struct {
		Reg#(Bit(32)) pc;
		Instr instr;
	} IfId;
		
	typedef struct {
	} IdEx;
		
	typedef struct {
	} ExMem;
		
	typedef struct {
	} MemWb;

endpackage
